// Create Date:    05/24/17
// Engineer(s):	   Triet Bach, Jim Lee, Aaron Yang
// Module Name:    Convert_Neg

module Conv_Neg (
   input [7:0] in,   
   output logic [7:0] out
   ); 

   assign out = -in;

endmodule 
